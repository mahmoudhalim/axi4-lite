package axi_lite_pkg;
    

typedef enum logic {IDLE, RADDR, RDATA, WADDR, WDATA, BRESP} state_e;

endpackage
